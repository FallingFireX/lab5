module circuit_b(
    input A, B, C, D, 
    output Y
);

   assign Y = //equation here

endmodule
